-- mips 32_bit single_cycle_processor
library ieee;
use ieee.std_logic_1164.all;
entity mips is  -- mips 32_bit single_cycle_processor  
    port(
        clk,rst : std_logic
    );
end entity;

architecture rtl of mips32_single_cycle is

end architecture;